case(i_coeff)
	0: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 10; end
			1: begin sign = 0; exp = 12; end
			2: begin sign = 0; exp = 14; end
		endcase
	end
	1: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 10; end
			1: begin sign = 1; exp = 14; end
		endcase
	end
	2: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 10; end
			1: begin sign = 0; exp = 13; end
			2: begin sign = 0; exp = 14; end
		endcase
	end
	3: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 10; end
			1: begin sign = 0; exp = 11; end
			2: begin sign = 0; exp = 14; end
		endcase
	end
	4: begin
		last = 1;
		case(i_term)
			0: begin sign = 0; exp = 9; end
		endcase
	end
	5: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 9; end
			1: begin sign = 0; exp = 11; end
		endcase
	end
	6: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 9; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 14; end
		endcase
	end
	7: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 1; exp = 11; end
		endcase
	end
	8: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 9; end
			1: begin sign = 0; exp = 11; end
			2: begin sign = 0; exp = 13; end
			3: begin sign = 0; exp = 14; end
		endcase
	end
	9: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 0; exp = 13; end
		endcase
	end
	10: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 0; exp = 11; end
			2: begin sign = 0; exp = 13; end
		endcase
	end
	11: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 13; end
		endcase
	end
	12: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 0; exp = 13; end
		endcase
	end
	13: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 8; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 12; end
		endcase
	end
	14: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 1; exp = 10; end
			2: begin sign = 1; exp = 13; end
		endcase
	end
	15: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 1; exp = 14; end
		endcase
	end
	16: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 0; exp = 10; end
		endcase
	end
	17: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 12; end
			3: begin sign = 0; exp = 13; end
		endcase
	end
	18: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 12; end
			3: begin sign = 0; exp = 13; end
		endcase
	end
	19: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 1; exp = 11; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	20: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 7; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 0; exp = 14; end
		endcase
	end
	21: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 1; exp = 9; end
			2: begin sign = 1; exp = 12; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	22: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 1; exp = 10; end
			2: begin sign = 1; exp = 12; end
		endcase
	end
	23: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 1; exp = 11; end
			2: begin sign = 1; exp = 13; end
		endcase
	end
	24: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 14; end
		endcase
	end
	25: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	26: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 1; exp = 11; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	27: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 0; exp = 14; end
		endcase
	end
	28: begin
		last = 5;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 0; exp = 9; end
			3: begin sign = 1; exp = 12; end
			4: begin sign = 1; exp = 14; end
		endcase
	end
	29: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 7; end
			2: begin sign = 1; exp = 10; end
			3: begin sign = 1; exp = 13; end
		endcase
	end
	30: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 7; end
			2: begin sign = 0; exp = 13; end
		endcase
	end
	31: begin
		last = 5;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 7; end
			2: begin sign = 0; exp = 10; end
			3: begin sign = 0; exp = 11; end
			4: begin sign = 0; exp = 13; end
		endcase
	end
	32: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 7; end
			2: begin sign = 0; exp = 10; end
			3: begin sign = 0; exp = 14; end
		endcase
	end
	33: begin
		last = 5;
		case(i_term)
			0: begin sign = 0; exp = 6; end
			1: begin sign = 0; exp = 7; end
			2: begin sign = 0; exp = 9; end
			3: begin sign = 0; exp = 11; end
			4: begin sign = 0; exp = 13; end
		endcase
	end
	34: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 8; end
			2: begin sign = 1; exp = 13; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	35: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 9; end
			2: begin sign = 1; exp = 10; end
			3: begin sign = 1; exp = 12; end
		endcase
	end
	36: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 9; end
			2: begin sign = 1; exp = 11; end
			3: begin sign = 0; exp = 14; end
		endcase
	end
	37: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 9; end
			2: begin sign = 0; exp = 12; end
		endcase
	end
	38: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 10; end
			2: begin sign = 1; exp = 13; end
		endcase
	end
	39: begin
		last = 2;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 1; exp = 12; end
		endcase
	end
	40: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 0; exp = 13; end
		endcase
	end
	41: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 10; end
			2: begin sign = 0; exp = 12; end
			3: begin sign = 0; exp = 13; end
		endcase
	end
	42: begin
		last = 3;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 1; exp = 13; end
		endcase
	end
	43: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 11; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	44: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 10; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	45: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 1; exp = 11; end
			3: begin sign = 1; exp = 13; end
		endcase
	end
	46: begin
		last = 4;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 8; end
			2: begin sign = 1; exp = 12; end
			3: begin sign = 1; exp = 14; end
		endcase
	end
	47: begin
		last = 5;
		case(i_term)
			0: begin sign = 0; exp = 5; end
			1: begin sign = 0; exp = 9; end
			2: begin sign = 0; exp = 10; end
			3: begin sign = 0; exp = 12; end
			4: begin sign = 0; exp = 14; end
		endcase
	end
endcase
